/// Display 4-bit binary to 2 led 7 doan

module part2(SW, HEX1, HEX0);
	input [3:0] SW;
	output [6:0] HEX1, HEX0;
	wire [0:0] s;
	wire [2:0] outA;
	wire [3:0] in1, in0;
	comparator compare(SW[3:0], s);
	circuitA circuit(SW[2:0], outA);
	assign in1 = (s ==1'b1) ? 4'b0001 : 4'b0000;
	assign in0 = (s == 1'b0) ? SW : outA;
	led_7seg hex1(in1, HEX1);
	led_7seg hex0(in0, HEX0);
endmodule
	

module comparator(SW, Z);
	input [3:0] SW;
	output [0:0] Z;
	assign Z = (SW == 4'b1010) ? 1:
			   (SW == 4'b1011) ? 1:
			   (SW == 4'b1100) ? 1:
			   (SW == 4'b1101) ? 1:
			   (SW == 4'b1110) ? 1:
			   (SW == 4'b1111) ? 1: 0;
endmodule

module circuitA(SW2_0, A);
	input [2:0] SW2_0;
	output [3:0] A;
	assign A = (SW2_0 == 3'b010) ? 4'b0000:
			   (SW2_0 == 3'b011) ? 4'b0001:
			   (SW2_0 == 3'b100) ? 4'b0010:
			   (SW2_0 == 3'b101) ? 4'b0011:
			   (SW2_0 == 3'b100) ? 4'b0100:
			   (SW2_0 == 3'b111) ? 4'b0101: 4'b1111;
endmodule

module led_7seg(in, Display);
	input [3:0] in;
	output [6:0] Display;
	assign Display = (in == 4'b0000) ? 7'b100_0000:
					 (in == 4'b0001) ? 7'b111_1001:
					 (in == 4'b0010) ? 7'b010_0100:
					 (in == 4'b0011) ? 7'b011_0000:
					 (in == 4'b0100) ? 7'b001_1001:
					 (in == 4'b0101) ? 7'b001_0010:
					 (in == 4'b0110) ? 7'b000_0010:
					 (in == 4'b0111) ? 7'b111_1000:
					 (in == 4'b1000) ? 7'b000_0000:
					 (in == 4'b1001) ? 7'b001_0000: 7'b111_1111;
endmodule

					 
	
