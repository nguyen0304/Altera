/// divide clock from 50MHz to 1Hz

module part3(Clk, Clk2);
	input Clk;
	output reg Clk2;
	
endmodule